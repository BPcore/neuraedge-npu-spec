// plusargs_router_stress.svh
`ifndef PLUSARGS_ROUTER_STRESS_SVH
`define PLUSARGS_ROUTER_STRESS_SVH
// +SEED=<n>          : RNG seed
// +INJECT_RATE=<n>   : average injection rate (packets/cycle * 1000)
// +BUILD_ONLY        : CI helper flag - build only
`endif // PLUSARGS_ROUTER_STRESS_SVH
