// uvm_traffic_seq.sv - example sequences for traffic/DVFS/sparsity
// Placeholders for sequence code that will drive CSR writes and traffic patterns.

// TODO: Implement sequence classes using your project's UVM base and CSR bus spec.

// Example pseudo-sequence:
// - write CSR util target to 0..100% in steps
// - inject traffic sequence with multi-destination masks
// - toggle sparsity modes and observe telemetry

// This file is a scaffold to be implemented when adopting a UVM flow.
