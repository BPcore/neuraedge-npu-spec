// Dummy property file for noc_router formal verification
// Add your SystemVerilog assertions here
module noc_router_props();
// ...property definitions...
endmodule
