// plusargs_dvfs_energy_convergence.svh
// Centralized plusargs / defaults for dvfs_energy_convergence_tb
`ifndef PLUSARGS_DVFS_ENERGY_CONVERGENCE_SVH
`define PLUSARGS_DVFS_ENERGY_CONVERGENCE_SVH
// Available plusargs (examples):
// +SEED=<n>           : RNG seed for randomized stimulus
// +SAMPLE_CYCLES=<n>  : number of energy sampling cycles (default 1000)
// +FORCE_UTIL=<pct>   : force a utilization value (0-100) for deterministic runs
// +BUILD_ONLY         : CI helper flag - build only, do not run long sim

`endif // PLUSARGS_DVFS_ENERGY_CONVERGENCE_SVH
