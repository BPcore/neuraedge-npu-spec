#
# NeuraEdge NPU - Final LEF Abstract Library for P&R Handoff  
# Phase 4 Week 4 Day 5: Freeze & Handoff
# Generated: August 14, 2025
# Status: FROZEN - Manufacturing Ready
#

################################################################################
# LEF HEADER AND TECHNOLOGY INFORMATION
################################################################################

VERSION 5.8 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

################################################################################
# TECHNOLOGY DEFINITION - TSMC 65nm GP
################################################################################

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.0 ;
  WIDTH 0.09 ;
  SPACING 0.09 ;
  RESISTANCE RPERSQ 0.38 ;
  CAPACITANCE CPERSQDIST 0.000207 ;
  THICKNESS 0.13 ;
  MINWIDTH 0.09 ;
  MAXWIDTH 2.0 ;
END M1

LAYER M2  
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.0 ;
  WIDTH 0.10 ;
  SPACING 0.10 ;
  RESISTANCE RPERSQ 0.38 ;
  CAPACITANCE CPERSQDIST 0.000164 ;
  THICKNESS 0.14 ;
  MINWIDTH 0.10 ;
  MAXWIDTH 2.0 ;
END M2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.0 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.27 ;
  CAPACITANCE CPERSQDIST 0.000133 ;
  THICKNESS 0.28 ;
  MINWIDTH 0.14 ;
  MAXWIDTH 4.0 ;
END M3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 2.0 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  RESISTANCE RPERSQ 0.27 ;
  CAPACITANCE CPERSQDIST 0.000133 ;
  THICKNESS 0.28 ;
  MINWIDTH 0.14 ;
  MAXWIDTH 4.0 ;
END M4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4.0 ;
  WIDTH 0.28 ;
  SPACING 0.28 ;
  RESISTANCE RPERSQ 0.19 ;
  CAPACITANCE CPERSQDIST 0.000108 ;
  THICKNESS 0.42 ;
  MINWIDTH 0.28 ;
  MAXWIDTH 8.0 ;
END M5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.0 ;
  WIDTH 0.28 ;
  SPACING 0.28 ;
  RESISTANCE RPERSQ 0.19 ;
  CAPACITANCE CPERSQDIST 0.000108 ;
  THICKNESS 0.42 ;
  MINWIDTH 0.28 ;
  MAXWIDTH 8.0 ;
END M6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 8.0 ;
  WIDTH 0.56 ;
  SPACING 0.56 ;
  RESISTANCE RPERSQ 0.09 ;
  CAPACITANCE CPERSQDIST 0.000087 ;
  THICKNESS 0.84 ;
  MINWIDTH 0.56 ;
  MAXWIDTH 16.0 ;
END M7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 8.0 ;
  WIDTH 0.56 ;
  SPACING 0.56 ;
  RESISTANCE RPERSQ 0.09 ;
  CAPACITANCE CPERSQDIST 0.000087 ;
  THICKNESS 0.84 ;
  MINWIDTH 0.56 ;
  MAXWIDTH 16.0 ;
END M8

################################################################################
# VIA DEFINITIONS
################################################################################

VIA VIA1
  LAYER M1 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER VIA1 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M2 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  RESISTANCE 4.5 ;
END VIA1

VIA VIA2
  LAYER M2 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER VIA2 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER M3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  RESISTANCE 2.1 ;
END VIA2

VIA VIA3
  LAYER M3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER VIA3 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER M4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  RESISTANCE 2.1 ;
END VIA3

VIA VIA4
  LAYER M4 ;
    RECT -0.070 -0.070 0.070 0.070 ;
  LAYER VIA4 ;
    RECT -0.140 -0.140 0.140 0.140 ;
  LAYER M5 ;
    RECT -0.140 -0.140 0.140 0.140 ;
  RESISTANCE 1.2 ;
END VIA4

VIA VIA5
  LAYER M5 ;
    RECT -0.140 -0.140 0.140 0.140 ;
  LAYER VIA5 ;
    RECT -0.140 -0.140 0.140 0.140 ;
  LAYER M6 ;
    RECT -0.140 -0.140 0.140 0.140 ;
  RESISTANCE 1.2 ;
END VIA5

VIA VIA6
  LAYER M6 ;
    RECT -0.140 -0.140 0.140 0.140 ;
  LAYER VIA6 ;
    RECT -0.280 -0.280 0.280 0.280 ;
  LAYER M7 ;
    RECT -0.280 -0.280 0.280 0.280 ;
  RESISTANCE 0.6 ;
END VIA6

VIA VIA7
  LAYER M7 ;
    RECT -0.280 -0.280 0.280 0.280 ;
  LAYER VIA7 ;
    RECT -0.280 -0.280 0.280 0.280 ;
  LAYER M8 ;
    RECT -0.280 -0.280 0.280 0.280 ;
  RESISTANCE 0.6 ;
END VIA7

################################################################################
# NEURAEDGE TILE MACRO DEFINITION
################################################################################

MACRO neuraedge_tile
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 500.0 BY 500.0 ;
  SYMMETRY X Y ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.0 498.0 500.0 500.0 ;
      LAYER M6 ;
        RECT 498.0 0.0 500.0 500.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 0.0 0.0 500.0 2.0 ;
      LAYER M6 ;
        RECT 0.0 0.0 2.0 500.0 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M4 ;
        RECT 248.0 0.0 252.0 4.0 ;
    END
  END CLK

  PIN RESET_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.0 0.0 247.0 4.0 ;
    END
  END RESET_N

  # Data interface pins (128-bit wide)
  PIN DATA_IN[127:0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 10.0 0.0 490.0 4.0 ;
    END
  END DATA_IN[127:0]

  PIN DATA_OUT[127:0]  
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 10.0 496.0 490.0 500.0 ;
    END
  END DATA_OUT[127:0]

  # NoC interface pins
  PIN NOC_NORTH_VALID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 240.0 496.0 244.0 500.0 ;
    END
  END NOC_NORTH_VALID

  PIN NOC_SOUTH_VALID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 240.0 0.0 244.0 4.0 ;
    END
  END NOC_SOUTH_VALID

  PIN NOC_EAST_VALID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 496.0 240.0 500.0 244.0 ;
    END
  END NOC_EAST_VALID

  PIN NOC_WEST_VALID
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 240.0 4.0 244.0 ;
    END
  END NOC_WEST_VALID

  # Memory interface pins
  PIN MEM_ADDR[31:0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.0 10.0 500.0 50.0 ;
    END
  END MEM_ADDR[31:0]

  PIN MEM_DATA[255:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.0 60.0 500.0 200.0 ;
    END
  END MEM_DATA[255:0]

  PIN MEM_CTRL[7:0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.0 210.0 500.0 230.0 ;
    END
  END MEM_CTRL[7:0]

  # Power control pins
  PIN POWER_GATE_CTRL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0 480.0 4.0 484.0 ;
    END
  END POWER_GATE_CTRL

  # Test and debug pins  
  PIN SCAN_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0 10.0 4.0 12.0 ;
    END
  END SCAN_IN

  PIN SCAN_OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 496.0 10.0 500.0 12.0 ;
    END
  END SCAN_OUT

  PIN SCAN_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0 14.0 4.0 16.0 ;
    END
  END SCAN_EN

  # Thermal monitoring
  PIN TEMP_SENSOR
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M1 ;
        RECT 480.0 480.0 484.0 484.0 ;
    END
  END TEMP_SENSOR

  OBS
    LAYER M1 ;
      RECT 20.0 20.0 480.0 480.0 ;
    LAYER M2 ;
      RECT 20.0 20.0 480.0 480.0 ;
    LAYER M3 ;
      RECT 20.0 20.0 480.0 480.0 ;
    LAYER M4 ;
      RECT 20.0 20.0 480.0 480.0 ;
  END

END neuraedge_tile

################################################################################
# SRAM 1MB MACRO DEFINITION
################################################################################

MACRO sram_1mb
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 100.0 BY 100.0 ;
  SYMMETRY X Y ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 0.0 98.0 100.0 100.0 ;
      LAYER M7 ;
        RECT 98.0 0.0 100.0 100.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M7 ;
        RECT 0.0 0.0 100.0 2.0 ;
      LAYER M7 ;
        RECT 0.0 0.0 2.0 100.0 ;
    END
  END VSS

  PIN VDD_RET
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 2.0 2.0 98.0 4.0 ;
    END
  END VDD_RET

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M5 ;
        RECT 48.0 0.0 52.0 4.0 ;
    END
  END CLK

  PIN ADDR[19:0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 10.0 0.0 40.0 4.0 ;
    END
  END ADDR[19:0]

  PIN DATA_IN[255:0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0 10.0 4.0 90.0 ;
    END
  END DATA_IN[255:0]

  PIN DATA_OUT[255:0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 96.0 10.0 100.0 90.0 ;
    END
  END DATA_OUT[255:0]

  PIN WE[31:0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 60.0 0.0 90.0 4.0 ;
    END
  END WE[31:0]

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 54.0 0.0 58.0 4.0 ;
    END
  END OE

  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 42.0 0.0 46.0 4.0 ;
    END
  END CE

  PIN POWER_GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 0.0 48.0 4.0 52.0 ;
    END
  END POWER_GATE

  PIN RETENTION_CTRL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 96.0 48.0 100.0 52.0 ;
    END
  END RETENTION_CTRL

  PIN BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0 92.0 4.0 96.0 ;
    END
  END BIST_EN

  PIN BIST_DONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.0 92.0 100.0 96.0 ;
    END
  END BIST_DONE

  PIN BIST_PASS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.0 88.0 100.0 92.0 ;
    END
  END BIST_PASS

  OBS
    LAYER M1 ;
      RECT 10.0 10.0 90.0 90.0 ;
    LAYER M2 ;
      RECT 10.0 10.0 90.0 90.0 ;
    LAYER M3 ;
      RECT 10.0 10.0 90.0 90.0 ;
  END

END sram_1mb

################################################################################
# NOC HUB MACRO DEFINITION
################################################################################

MACRO noc_hub
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 50.0 BY 50.0 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.0 48.0 50.0 50.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 0.0 0.0 50.0 2.0 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M5 ;
        RECT 24.0 0.0 26.0 4.0 ;
    END
  END CLK

  # Tile interface ports (4x4 = 16 ports)
  PIN TILE_NORTH[15:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.0 46.0 45.0 50.0 ;
    END
  END TILE_NORTH[15:0]

  PIN TILE_SOUTH[15:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.0 0.0 45.0 4.0 ;
    END
  END TILE_SOUTH[15:0]

  PIN TILE_EAST[15:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 46.0 5.0 50.0 45.0 ;
    END
  END TILE_EAST[15:0]

  PIN TILE_WEST[15:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 5.0 4.0 45.0 ;
    END
  END TILE_WEST[15:0]

  # Memory interface ports
  PIN MEM_NORTH[63:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 10.0 40.0 40.0 46.0 ;
    END
  END MEM_NORTH[63:0]

  PIN MEM_SOUTH[63:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 10.0 4.0 40.0 10.0 ;
    END
  END MEM_SOUTH[63:0]

  # I/O interface ports  
  PIN IO_INTERFACE[31:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 20.0 20.0 30.0 30.0 ;
    END
  END IO_INTERFACE[31:0]

  OBS
    LAYER M1 ;
      RECT 5.0 5.0 45.0 45.0 ;
    LAYER M2 ;
      RECT 5.0 5.0 45.0 45.0 ;
  END

END noc_hub

################################################################################
# NOC ROUTER MACRO DEFINITION
################################################################################

MACRO noc_router
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 25.0 BY 25.0 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 0.0 23.0 25.0 25.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 0.0 0.0 25.0 2.0 ;
    END
  END VSS

  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M4 ;
        RECT 11.0 0.0 14.0 4.0 ;
    END
  END CLK

  PIN ROUTER_NORTH[31:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5.0 21.0 20.0 25.0 ;
    END
  END ROUTER_NORTH[31:0]

  PIN ROUTER_SOUTH[31:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 5.0 0.0 20.0 4.0 ;
    END
  END ROUTER_SOUTH[31:0]

  PIN ROUTER_EAST[31:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 21.0 5.0 25.0 20.0 ;
    END
  END ROUTER_EAST[31:0]

  PIN ROUTER_WEST[31:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0 5.0 4.0 20.0 ;
    END
  END ROUTER_WEST[31:0]

  OBS
    LAYER M1 ;
      RECT 2.0 2.0 23.0 23.0 ;
    LAYER M2 ;
      RECT 2.0 2.0 23.0 23.0 ;
  END

END noc_router

################################################################################
# I/O CONTROLLER MACRO DEFINITION  
################################################################################

MACRO io_controller
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 50.0 BY 25.0 ;

  PIN VDD_IO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 0.0 23.0 50.0 25.0 ;
    END
  END VDD_IO

  PIN VDD_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.0 21.0 50.0 23.0 ;
    END
  END VDD_CORE

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M7 ;
        RECT 0.0 0.0 50.0 2.0 ;
    END
  END VSS

  PIN CLK_IO
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M5 ;
        RECT 24.0 0.0 26.0 4.0 ;
    END
  END CLK_IO

  PIN IO_DATA[63:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 5.0 0.0 45.0 4.0 ;
    END
  END IO_DATA[63:0]

  PIN IO_CTRL[15:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 10.0 21.0 40.0 25.0 ;
    END
  END IO_CTRL[15:0]

  PIN CORE_INTERFACE[127:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0 10.0 4.0 15.0 ;
    END
  END CORE_INTERFACE[127:0]

  OBS
    LAYER M1 ;
      RECT 5.0 5.0 45.0 20.0 ;
    LAYER M2 ;
      RECT 5.0 5.0 45.0 20.0 ;
  END

END io_controller

################################################################################
# CLOCK BUFFER MACRO DEFINITIONS
################################################################################

MACRO clock_buffer_x16
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 10.0 BY 10.0 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0.0 8.0 10.0 10.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0.0 0.0 10.0 2.0 ;
    END
  END VSS

  PIN CLK_IN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 0.0 4.0 2.0 6.0 ;
    END
  END CLK_IN

  PIN CLK_OUT
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 8.0 4.0 10.0 6.0 ;
    END
  END CLK_OUT

  OBS
    LAYER M1 ;
      RECT 2.0 2.0 8.0 8.0 ;
  END

END clock_buffer_x16

MACRO clock_buffer_x8
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 8.0 BY 8.0 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0.0 6.0 8.0 8.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0.0 0.0 8.0 2.0 ;
    END
  END VSS

  PIN CLK_IN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 0.0 3.0 2.0 5.0 ;
    END
  END CLK_IN

  PIN CLK_OUT
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 6.0 3.0 8.0 5.0 ;
    END
  END CLK_OUT

  OBS
    LAYER M1 ;
      RECT 2.0 2.0 6.0 6.0 ;
  END

END clock_buffer_x8

################################################################################
# POWER MANAGEMENT MACRO DEFINITIONS
################################################################################

MACRO power_mgmt_unit
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 20.0 BY 20.0 ;

  PIN VDD_AON
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M7 ;
        RECT 0.0 18.0 20.0 20.0 ;
    END
  END VDD_AON

  PIN VDD_SWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 0.0 16.0 20.0 18.0 ;
    END
  END VDD_SWITCH

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M7 ;
        RECT 0.0 0.0 20.0 2.0 ;
    END
  END VSS

  PIN CLK_AON
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M5 ;
        RECT 9.0 0.0 11.0 4.0 ;
    END
  END CLK_AON

  PIN POWER_CTRL[7:0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0 8.0 4.0 12.0 ;
    END
  END POWER_CTRL[7:0]

  PIN POWER_STATUS[7:0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.0 8.0 20.0 12.0 ;
    END
  END POWER_STATUS[7:0]

  PIN VOLTAGE_MON[3:0]
    DIRECTION OUTPUT ;
    USE ANALOG ;
    PORT
      LAYER M3 ;
        RECT 8.0 16.0 12.0 20.0 ;
    END
  END VOLTAGE_MON[3:0]

  OBS
    LAYER M1 ;
      RECT 4.0 4.0 16.0 16.0 ;
    LAYER M2 ;
      RECT 4.0 4.0 16.0 16.0 ;
  END

END power_mgmt_unit

################################################################################
# DEBUG AND TEST MACRO DEFINITIONS
################################################################################

MACRO debug_ctrl
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 15.0 BY 15.0 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 0.0 13.0 15.0 15.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 0.0 0.0 15.0 2.0 ;
    END
  END VSS

  PIN DEBUG_CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M4 ;
        RECT 7.0 0.0 8.0 4.0 ;
    END
  END DEBUG_CLK

  PIN DEBUG_DATA[31:0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0 5.0 4.0 10.0 ;
    END
  END DEBUG_DATA[31:0]

  PIN DEBUG_CTRL[7:0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 11.0 5.0 15.0 7.0 ;
    END
  END DEBUG_CTRL[7:0]

  OBS
    LAYER M1 ;
      RECT 3.0 3.0 12.0 12.0 ;
  END

END debug_ctrl

MACRO jtag_ctrl
  CLASS BLOCK ;
  ORIGIN 0.0 0.0 ;
  SIZE 12.0 BY 12.0 ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0.0 10.0 12.0 12.0 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 0.0 0.0 12.0 2.0 ;
    END
  END VSS

  PIN TCK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M3 ;
        RECT 0.0 5.0 2.0 7.0 ;
    END
  END TCK

  PIN TDI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0 3.0 2.0 5.0 ;
    END
  END TDI

  PIN TDO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 10.0 5.0 12.0 7.0 ;
    END
  END TDO

  PIN TMS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0 7.0 2.0 9.0 ;
    END
  END TMS

  PIN TRST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0 9.0 2.0 10.0 ;
    END
  END TRST_N

  OBS
    LAYER M1 ;
      RECT 2.0 2.0 10.0 10.0 ;
  END

END jtag_ctrl

################################################################################
# SITE DEFINITIONS FOR STANDARD CELLS
################################################################################

SITE CoreSite
  CLASS CORE ;
  SIZE 0.6 BY 4.0 ;
END CoreSite

SITE IOSite
  CLASS PAD ;
  SIZE 100.0 BY 100.0 ;
END IOSite

SITE MemorySite
  CLASS BLOCK ;
  SIZE 100.0 BY 100.0 ;
END MemorySite

################################################################################
# DESIGN RULES
################################################################################

PROPERTYDEFINITIONS
  DESIGN FOREIGN STRING ;
  LAYER MANUFACTURINGGRID REAL ;
  LAYER MAXWIDTH REAL ;
  LAYER MINWIDTH REAL ;
  MACRO FOREIGN STRING ;
  PIN FOREIGN STRING ;
END PROPERTYDEFINITIONS

MANUFACTURINGGRID 0.005 ;

################################################################################
# LEF FILE CLOSURE
################################################################################

END LIBRARY
