`timescale 1ns/1ps
// Skeleton NoC random stress TB (to be completed): will drive random flits into mesh ends
module noc_random_stress_tb;
  initial begin
    $display("[NOC_RAND] Placeholder start");
    #20;
    $display("[NOC_RAND] Placeholder end");
    $finish;
  end
endmodule
