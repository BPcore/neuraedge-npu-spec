// uvm_csr_agent.sv - CSR agent scaffold (UVM)
// This is a skeleton to be expanded into full UVM driver/monitor/agent.

// NOTE: This file is intentionally minimal; implement UVM classes (uvm_driver, uvm_monitor, etc.) when using a UVM simulator.

// Placeholder package guard
`ifndef UVM_CSR_AGENT_SV
`define UVM_CSR_AGENT_SV

// ... UVM implementation goes here ...

`endif
