// sequences/uvm_csr_seq.sv
// Minimal UVM sequence scaffold: perform a few CSR reads/writes as a sanity sequence.

`ifndef UVM_CSR_SEQ_SV
`define UVM_CSR_SEQ_SV

// Sequence placeholder; expand for real UVM usage.

`endif
