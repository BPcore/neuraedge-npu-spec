// uvm_env.sv - minimal UVM environment scaffold
`ifndef UVM_ENV_SV
`define UVM_ENV_SV

// Minimal placeholder env - expand with real UVM components when targeting a UVM-capable simulator.
module uvm_env_svb;
  // Placeholder wrapper to hold UVM env files for source control and incremental implementation.
  // See README.md for guidance on next steps.
endmodule

`endif
