// Physical synthesis placeholder - base netlist not available
module neuraedge_top(); endmodule
