// File: rtl/top/neuraedge_top.sv
module neuraedge_top (
  input  logic        clk,
  input  logic        rst_n
  // TODO: add tile instantiations, NoC interconnect, external I/O ports
);

  // Stub: nothing yet, just a placeholder to satisfy lint
  // All actual ports and signals will be added in Week 3

endmodule
