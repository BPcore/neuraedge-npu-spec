// plusargs_mem_contention.svh
`ifndef PLUSARGS_MEM_CONTENTION_SVH
`define PLUSARGS_MEM_CONTENTION_SVH
// +SEED=<n>             : RNG seed
// +REQUESTS_PER_TILE=<n>: number of requests per tile in deterministic variants
// +QUEUE_DEPTH=<n>      : injector queue depth override
// +BUILD_ONLY           : CI helper flag - build only
`endif // PLUSARGS_MEM_CONTENTION_SVH
